`timescale 1ns / 1ps

module Data_codec(
	input r_enable,
	input [0:95] m_data,
	input [0:2] linesel,
	
	output reg linesel_en,
	output reg [0:31]red,
	output reg [0:31]red2,
	output send,
	output enable
    );


	integer i, u_i=0, u_f=2, a;
	reg[0:7]matrix_R[31:0];
	reg[0:7]data_c;
	reg [0:95] data_desp;
	
initial begin	
data_desp<= m_data;

	while(r_enable==1) begin
	linesel_en<=0;
	for (i=0;i<=31;i=i+1) begin
	
	a<=data_desp[0:2];
	data_desp<= data_desp<<3;
		//u_i<=u_i+2'd3;
		//u_f<=u_f+2'd3;
//		a<=m_data[u_i];
//		u_i<=u_i+2'd3;
//		u_f<=u_f+2'd3;
		
		case(a)
			0: data_c=8'd128;
			1: data_c=8'd192;
			2: data_c=8'd224;
			3: data_c=8'd240;
			4: data_c=8'd248;
			5: data_c=8'd252;
			6: data_c=8'd254;
			7: data_c=8'd255;
			default: data_c=8'd255;
		endcase
	
		matrix_R[i]=data_c;
	
	end //for
	end //while
	
	linesel_en<=1;
	
	while(linesel==0) begin
		red=matrix_R[0][0:31];
		red2=matrix_R[7][0:31];
	end
	while(linesel==1) begin
		red=matrix_R[1][0:31];
		red2=matrix_R[6][0:31];
	end
	while(linesel==2) begin
		red=matrix_R[2][0:31];
		red2=matrix_R[5][0:31];
	end
	while(linesel==3) begin
		red=matrix_R[3][0:31];
		red2=matrix_R[4][0:31];
	end
	while(linesel==4) begin
		red=matrix_R[4][0:31];
		red2=matrix_R[3][0:31];
	end
	while(linesel==5) begin
		red=matrix_R[5][0:31];
		red2=matrix_R[2][0:31];
	end
	while(linesel==6) begin
		red=matrix_R[6][0:31];
		red2=matrix_R[1][0:31];
	end
	while(linesel==7) begin
		red=matrix_R[7][0:31];
		red2=matrix_R[0][0:31];
	end
end

endmodule
